LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.std_logic_signed.all;

ENTITY OU IS

PORT ( 
X, Y : IN STD_LOGIC_VECTOR(7 DOWNTO 0) ;
S : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) 
 ) ;
END OU ;
ARCHITECTURE logica OF OU IS

BEGIN

S <= X OR Y;


END logica ;